5�d d         d    ��  CprobeN  ����b  ����[  ����q  ����  A     ��  CpinX  ����X  ����0 0 A[  ����          �U  "���i  ���b  4���x  "���  B     �_  ���_  ���0 0 Bb  4���          �g  x���{  X���t  �����  x���  C     �q  X���q  f���0 0 Ct  ����          �� 
 CDflipflop�  �����  ?���                       ��  e����  e���0 0                  ��  }����  }���Z Z                  ��  �����  ����1 1                  ��  ?����  M���1 1                   ��  }����  }���0 0                  ��  e����  e���1 1                  	��  ���   ����                       ��  �����  ����0 0                  ��  �����  ����0 0                  ��  ����  ����1 1                  ��  �����  ����1 1                   �   �����  ����0 0                  �   �����  ����1 1                  	��  n���  
���                       ��  0����  0���0 0                  ��  H����  H���X X                  ��  n����  `���1 1                  ��  
����  ���1 1                   �  H����  H���0 0                  �  0����  0���1 1                  ��  CswitchM  ����Y  ����c  �����  ���� Clock    �Y  ����Y  ����1 }                  �M  ����M  ����0 ��                  �S  ����S  ����0 0 Clockc  ����        ��  ����.  ����  ����6  ���� PreA    �.  ����   ����1 _                  �.  ����   ����0 `                   ��  ����  ����1 0 PreA  ����        ��  ���)  ���  0���1  ��� PreB    �)  ���  ���1 b                  �)  ���  ���0 c                   ��  ���  ���1 0 PreB  0���        ��  o���.  c���  ����6  o��� PreC    �.  c���   c���1 f                  �.  o���   o���0 g                   ��  i���  i���1 0 PreC  ����        �O  ����[  ����e  �����  ���� CirALL    �O  ����O  ����1 [                  �[  ����[  ����0 \                   �U  ����U  ����1 0 CirALLe  ����        �� 	 Cinverterf  �����  ����                       �f  ����t  ����1 1                   ��  �����  ����0 0                  ��  Cnand2�   ����F  ����                       ��   ����	  ����0 0                  ��   ����	  ����1 1                   �E  ����7  ����1 1                  8�k  Z����  6���                       �k  N���y  N���X X                  �k  B���y  B���X X                   ��  H����  H���X X                  4��   ~���7  Z���                       ��   l���  l���Z Z                   �7  l���)  l���X X                  4��   S���:  /���                       ��   A���
  A���Z Z                   �:  A���,  A���X X                   ��  Cnet0  ��  CsegmentS  ����S  +���I�S  ����S  ����I�S  +����  +���I��  0����  +���I��  0����  0���I�S  e����  e���I�S  ����S  e���I��  e����  e���I�S  �����  ����I�S  e���S  ����I��  �����  ����     # G�0  I�X  ����X  }���I��  }���X  }���I��  }����  }���I�X  ����X  ����    G�0  I�_  ���_  ����I�   ����_  ����I�   ����   ����I�_  ���_  ���    G�0 
 I�q  X���q  H���I�  H���q  H���I�  H���  H���I�q  X���q  X���I�  H���  H���I�  ����  H���I��   �����   ����I��   �����   ����I��   ����  ����I��   �����   ����  :   G�1  I��  �����  ����I��  �����  ����I��  �����  ����I��  �����  ����   ' G�1  I��  ����  ���I��  ����  ���I��  ����  ���I��  ����  ���   + G�1  I��  n����  i���I��  i����  i���I��  i����  i���I��  n����  n���   / G�1  I��  
����  ����I�=  �����  ����I�U  ����U  ����I��  
����  
���I�U  ����=  ����I�=  ����=  ?���I��  ?���=  ?���I��  ?����  ?���I�=  �����  ����I�=  ����=  ����I��  �����  ����     3 G�0  I��  �����  ����I��  �����  ����I��  �����  ����I��  �����  ����   7 G�1  I�   ����   ����I�  ����   ����I�  ����  ����I��   �����   ����I��   �����   ����I�  �����   ���� ;   G�1  I�f  ����f  ����I�E  ����f  ����I�E  ����E  ����I�f  ����f  ���� 6  < G�X  I��  H����  H���I��  H����  H���I��  H����  H���   @ G�X  I�k  B���k  B���I�;  A���:  A���I�:  A���:  A���I�;  A���;  8���I�;  B���;  A���I�k  B���;  B��� ?  F G�X  I�F  l���F  l���I�k  N���k  N���I�F  l���7  l���I�F  N���F  l���I�7  l���7  l���I�k  N���F  N��� >  C   joshua