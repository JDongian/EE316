5�d d         d    ��  Cprobe�  �����  �����  �����  ����  A     ��  Cpin�  �����  ����0 0 A�  ����          ��   ����   ����  2����   ���  B     ��   ����  ���0 0 B�   ���          ��  v����  V����  �����  v���  C     ��  V����  d���0 0 C�  V���          �� 
 CDflipflop  ����X  =���                       �  c���"  c���0 0                  �  {���"  {���Z Z                  �6  ����6  ����0 0                  �6  =���6  K���0 0                   �X  {���J  {���0 0                  �X  c���J  c���1 1                  	�  	���\  ����                       �  ����&  ����0 0                  �  ����&  ����Z Z                  �:  	���:  ����0 0                  �:  ����:  ����0 0                   �\  ����N  ����0 0                  �\  ����N  ����1 1                  	�  l���a  ���                       �  .���+  .���0 0                  �  F���+  F���Z Z                  �?  l���?  ^���0 0                  �?  ���?  ���0 0                   �a  F���S  F���0 0                  �a  .���S  .���1 1                  ��  Cswitch�   �����   �����   �����   ���� Clock    ��   �����   ����1 }                  ��   �����   ����0 ��                  ��   �����   ����0 0 Clock�   ����        �Z  �����  ����g  �����  ���� PreA    ��  ����|  ����1 _                  ��  ����|  ����0 `                   �Z  ����h  ����0 0 PreAB  ����        �U  ����  ���b  .����  ��� PreB    ��  ���w  ���1 b                  ��  ���w  ���0 c                   �U  ���c  ���0 0 PreB=  #���        �Z  m����  a���g  ����  m��� PreC    ��  a���|  a���1 f                  ��  m���|  m���0 g                   �Z  g���h  g���0 0 PreCB  t���        ��  �����  �����  �����  ���� CirALL    ��  �����  ����1 [                  ��  �����  ����0 \                   ��  �����  ����0 0 CirALL�  ����         ��  Cnet0  ��  Csegment�   �����   )���6��   �����   ����6��   )���  )���6�  .���  )���6�  .���  .���6��   c���  c���6��   �����   c���6�  c���  c���6��   ����  ����6��   c����   ����6�  ����  ����     # 4�0  6��  �����  {���6�X  {����  {���6�X  {���X  {���6��  �����  ����    4�0  6��   ����  ����6�\  �����  ����6�\  ����\  ����6��   ����   ���    4�0  6��  V����  F���6�a  F����  F���6�a  F���a  F���6��  V����  V���    4�0  6�6  ����6  ����6�Z  ����6  ����6�Z  ����Z  ����6�6  ����6  ����   ' 4�0  6�:  	���:  ���6�U  ���:  ���6�U  ���U  ���6�:  	���:  	���   + 4�0  6�?  l���?  g���6�Z  g���?  g���6�Z  g���Z  g���6�?  l���?  l���   / 4�0  6�?  ���?  ����6��  ����?  ����6��  �����  ����6�?  ���?  ���6��  �����  ����6��  �����  =���6�6  =����  =���6�6  =���6  =���6��  ����:  ����6��  �����  ����6�:  ����:  ����     3   joshua