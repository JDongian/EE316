5�         d    ��  Cprobef  ����  ����j  �����  ����  Q1     ��  Cpins  ����s  ����0 0 Q1j  ����          �n  �����  ����n  ����  ����  Q2     �{  ����{  ����0 0 Q2n  ���          ��  '����  �����  <����  %���  Q3     ��  �����  ���1 1 Q3�  <���          �� 
 CDflipflop�  �����  6���                       ��  f����  f���0 0                  ��  �����  ����0 0                  ��  �����  ����1 1                  ��  6����  G���1 1                   ��  �����  ����0 0                  ��  f����  f���1 1                  	��  ����  u���                       ��  �����  ����0 0                  ��  �����  ����1 1                  ��  �����  ����1 1                  ��  u����  ����1 1                   �  �����  ����0 0                  �  �����  ����1 1                  	��  -���	  ����                       ��  �����  ����0 0                  ��  �����  ����0 0                  ��  -����  ���1 1                  ��  �����  ����1 1                   �	  �����  ����1 1                  �	  �����  ����0 0                  ��  Cswitch!  ����0  ����=  ����k  ���� clk    �0  ����0  ����1 }                  �!  ����!  ����0 ��                  �(  ����(  ����0 0 clk=  ����        ��  ����9  ����                      �9  ����(  ����1 _                  �9  ����(  ����0 `                   ��  ����  ����1 0                  ��  ���7  ����                      �7  ����%  ����1 b                  �7  ���%  ���0 c                   ��  ���  ���1 0                  �   4���=  %���                      �=  %���,  %���1 f                  �=  4���,  4���0 g                   �   -���  -���1 0                  �H  a���W  %���e  E����  .��� rst    �H  %���H  6���1 [                  �W  %���W  6���0 \                   �P  a���P  P���1 0 rste  E���        �   ����K   ����    ����<   ���� x     �   ����!   ����1                    �   ����!   ����0                     �K   ����:   ����0 0 x    ����        �#  ����<  ����4  ����P  ����  Z     �0  ����0  ����1 1 Z4  ����          ��  Cnor3@  �����  ����                       �@  ����X  ����0 0                  �@  ����Z  ����0 0                  �@  ����X  ����0 0                   ��  �����  ����1 1                  ��  Cnand2�  ����  ����                       ��  �����  ����1 1                  ��  �����  ����0 0                   �  ����   ����1 1                  �� 	 Cinverter�   �����   ����                       ��   �����   ����0 0                   ��   �����   ����1 1                  @�D  ����  ����                       �D  ���U  ���1 1                  �D  ����U  ����1 1                   ��  �����  ����0 0                  @��   ����   ����                       ��   �����   ����0 0                  ��   �����   ����1 1                   ��   �����   ����1 1                  ��  Cnand3�   M����    ���                       ��   F����   F���1 1                  ��   7����   7���1 1                  ��   '����   '���0 0                   ��   7����   7���1 1                  @�,  4����  ���                       �,  %���=  %���0 0                  �,  ���=  ���0 0                   ��  ���w  ���1 1                  @�+  �����  ����                       �+  ����<  ����1 1                  �+  ����<  ����1 1                   ��  ����v  ����0 0                   ��  Cnet0 
 ��  Csegment(  ����(  ����a�(  ����(  ����a��  �����  ����a�(  f����  f���a��  f����  f���a�(  �����  ����a�(  f���(  ����a��  �����  ����a�(  �����  ����a�(  ����(  f���     # _�0 	 a�  ����s  ����a��  �����  ����a�s  ����s  ����a��  ����  ����a�  ����  ���a�  ���  ���a�  ���  ����a�@  ����  ����a�@  ����@  ����  <   _�0  a�{  ����{  ����a�{  ����{  ����a�  ����  ����a�  ����{  ����a�  ����  ����a�  ����  Y���a��   Y���  Y���a��   �����   ����a��  �����   ����a��  �����  ����a��   �����   Y���a�@  ����@  ����a��   ����@  ����   =   _�1  a��  �����  ����a��  �����  ����a��  �����  ����a��  �����  ����   ' _�1  a��  �����  ���a��  ����  ���a��  ����  ���a��  �����  ����   + _�1  a�   -���   -���a��  -����  -���a�   -����  -���   / _�1  a��  �����  ����a�P  �����  ����a�P  a���P  a���a��  �����  ����a�P  u���P  6���a��  6���P  6���a��  6����  6���a�P  u����  u���a�P  ����P  u���a��  u����  u���a�P  a���P  ����     3 _�0  a�@  ����@  ����a�  ����@  ����a�  ���  s���a�	  s���  s���a�  s���  ���a�,  ���  ���a�	  ����	  s���a�	  ����	  ����a�  ����  ���a�  ����   ���a��   '����   ���a��   '����   '���a�,  ���,  ��� > U Y   _�1  a��  �����  ����a��  �����  ����a��  �����  ����   ? _�Z       _�1  a�0  ����0  ����a�  ����  ����a�0  ����0  ����a�  ����0  ���� 9  D _�0  a�k   �����   ����a��   %����   ����a�K   ����K   ����a��   �����   ����a��   %����   ����a��   �����   ����a��   %���,  %���a�K   ����k   ����a�k   ����k   ����a��   ����k   ����a��   �����   ����a�,  %���,  %��� G N X  7 _�Z  a�  ����  ����    _�Z       _�1  a��   �����   ����a�D  ����D  ����a��   ����D  ���� K  P _�1  a��   ����   7���a�D  ���D  ���a��   ���D  ���a��   7����   7���a��   7����   7��� J  V _�0  a��  �����  ����a��  �����  ����a��  �����  ����   L _�1  a�  ����  e���a�  ����  ����a�  e���~   e���a�~   7���~   e���a��   7����   7���a�~   7����   7��� T   _�1  a��  f���  f���a�  *���  f���a��  f����  f���a�  *���n   *���a�n   F���n   *���a��   F����   F���a�n   F����   F��� S   _�0  a��  �����  ����a��  �����  ����a��  �����  ����a��  �����  ���� C  ^ _�Z       _�1  a�0  ����0  ����a��  �����  ����a��  �����  ����a��  ����  ����a�  ����	  ����a�  ����  c���a�  c���  c���a�  ����  c���a�  ����z   ����a�z   ����z   ����a�z   �����   ����a��   �����   ����a�	  ����	  ����a�  ����  c���a�  ����+  ���� ]  O   _�1  a��   ����+  ����a��   �����   �����  \  H _�1  a��  ����  ���a��  ����  ���a��  �����  ����a��  �����  ����a��  �����  ��� B  Z   joshua