5�d d         d    ��  CprobeN  ����b  ����[  ����q  ����  A     ��  CpinX  ����X  ����0 0 A[  ����          �U  "���i  ���b  4���x  "���  B     �_  ���_  ���0 0 Bb  4���          �g  x���{  X���t  �����  x���  C     �q  X���q  f���0 0 Ct  ����          �� 
 CDflipflop�  �����  ?���                       ��  e����  e���0 0                  ��  }����  }���Z Z                  ��  �����  ����1 1                  ��  ?����  M���1 1                   ��  }����  }���0 0                  ��  e����  e���1 1                  	��  ���   ����                       ��  �����  ����0 0                  ��  �����  ����0 0                  ��  ����  ����1 1                  ��  �����  ����1 1                   �   �����  ����0 0                  �   �����  ����1 1                  	��  n���  
���                       ��  0����  0���0 0                  ��  H����  H���1 1                  ��  n����  `���1 1                  ��  
����  ���1 1                   �  H����  H���0 0                  �  0����  0���1 1                  ��  CswitchM  ����Y  ����c  �����  ���� Clock    �Y  ����Y  ����1 }                  �M  ����M  ����0 ��                  �S  ����S  ����0 0 Clockc  ����        ��  ����.  ����  ����6  ���� PreA    �.  ����   ����1 _                  �.  ����   ����0 `                   ��  ����  ����1 0 PreA  ����        ��  ���)  ���  %���1  ��� PreB    �)  ���  ���1 b                  �)  ���  ���0 c                   ��  ���  ���1 0 PreB  %���        ��  s���.  g���  ����6  s��� PreC    �.  g���   g���1 f                  �.  s���   s���0 g                   ��  m���  m���1 0 PreC  ����        �O  ����[  ����e  �����  ���� CirALL    �O  ����O  ����1 [                  �[  ����[  ����0 \                   �U  ����U  ����1 0 CirALLe  ����        �� 	 Cinverterf  �����  ����                       �f  ����t  ����1 1                   ��  �����  ����0 0                  ��  Cnand2�   ����F  ����                       ��   ����	  ����0 0                  ��   ����	  ����1 1                   �E  ����7  ����1 1                  8�k  Z����  6���                       �k  N���y  N���0 0                  �k  B���y  B���0 0                   ��  H����  H���1 1                  4��   ~���:  Z���                       ��   l���
  l���1 1                   �:  l���,  l���0 0                  4��   T���:  0���                       ��   B���
  B���1 1                   �:  B���,  B���0 0                  8��   ~����   Z���                       ��   r����   r���0 0                  ��   f����   f���1 1                   ��   l����   l���1 1                  8��   S����   /���                       ��   G����   G���0 0                  ��   ;����   ;���1 1                   ��   A����   A���1 1                   ��  Cnet0 
 ��  CsegmentS  0���S  ����Q�S  ����S  ����Q��  0����  0���Q�S  e����  e���Q�S  ����S  e���Q��  e����  e���Q�S  �����  ����Q�S  e���S  ����Q��  �����  ����Q��  0���S  0���     # O�0 
 Q�X  ����X  }���Q�  }���X  }���Q��  }����  }���Q�X  ����X  ����Q��  }���  }���Q�  }���  $���Q�c   $���  $���Q�c   $���c   G���Q��   G���c   G���Q��   G����   G���  L   O�0 
 Q�_  ���_  ����Q�  ����_  ����Q�   ����   ����Q�_  ���_  ���Q�   ����  ����Q�  ����  ����Q��   ����  ����Q��   �����   r���Q��   r����   r���Q��   r����   r���  H   O�0 
 Q�q  X���q  H���Q�  H���q  H���Q�  H���  H���Q�q  X���q  X���Q�  H���  ����Q��   �����   ����Q��   �����   ����Q��   ����  ����Q��   �����   ����Q�  H���  H���  :   O�1  Q��  �����  ����Q��  �����  ����Q��  �����  ����Q��  �����  ����   ' O�1  Q��  ����  ���Q��  ����  ���Q��  ����  ���Q��  ����  ���Q��  ����  ���   + O�1  Q��  m����  m���Q��  n����  n���Q��  m����  n���Q��  n����  n���   / O�1  Q��  ����=  ����Q�U  ����U  ����Q��  
����  
���Q�U  ����=  ����Q�=  ����=  ?���Q��  ?���=  ?���Q��  ?����  ?���Q�=  �����  ����Q�=  ����=  ����Q��  �����  ����Q��  
����  ����     3 O�0  Q��  �����  ����Q��  �����  ����Q��  �����  ����Q��  �����  ����   7 O�1  Q�   ����   ����Q�  ����   ����Q�  ����  ����Q��   �����   ����Q��   �����   ����Q�  �����   ����Q��   ����o   ����Q�o   <���o   ����Q��   <����   ;���Q��   ;����   ;���Q�o   <����   <��� ; M   O�1  Q�f  ����f  ����Q�E  ����f  ����Q�E  ����E  ����Q�f  ����f  ���� 6  < O�1  Q��  H����  H���Q��  H����  H���Q��  H����  H���   @ O�Z       O�0  Q�:  B���k  B���Q�k  B���k  B���Q�:  B���:  B��� ?  F O�0  Q�:  l���:  N���Q�k  N���:  N���Q�k  N���k  N���Q�:  l���:  l��� >  C O�1  Q��   l����   l���Q��   l����   l���Q��   l����   l��� B  J O�1  Q��   B����   A���Q��   A����   A���Q��   A����   A���Q��   B����   B��� E  N O�1  Q�  0���  0���Q�  ����}   ����Q�}   f���}   ����Q��   f����   f���Q�  0���  ����Q�}   f����   f���Q�  0���  0��� I     joshua