5�d d        d    ��  CprobeV  ����j  ����c  ����  ����  Q1     ��  Cpin`  ����`  ����0 0 Q1c  ����          �]  ���q  ����j   ����  ���  Q2     �g  ����g  ����0 0 Q2j   ���          �r  e����  E���  w����  e���  Q3     �|  E���|  S���1 1 Q3  w���          �� 
 CDflipflop�  ����  +���                       ��  Q����  Q���1 1                  ��  i����  i���0 0                  ��  �����  ����1 1                  ��  +����  9���1 1                   �  i����  i���0 0                  �  Q����  Q���1 1                  	��  ����  ����                       ��  �����  ����1 1                  ��  �����  ����0 0                  ��  �����  ����1 1                  ��  �����  ����1 1                   �  �����  ����0 0                  �  �����  ����1 1                  	��  Z���  ����                       ��  ����  ���1 1                  ��  4����  4���1 1                  ��  Z����  L���1 1                  ��  �����  ���1 1                   �  4����  4���1 1                  �  ����  ���0 0                  ��  CswitchU  ����a  ����k  �����  ���� Clock    �a  ����a  ����1 }                  �U  ����U  ����0 ��                  �[  ����[  ����1 0 Clockk  ����        �  ����6  ����  ����>  ���� PreA    �6  ����(  ����1 _                  �6  ����(  ����0 `                   �  ����  ����1 0 PreA  ����        �  
���1  ����  ���9  
��� PreB    �1  ����#  ����1 b                  �1  
���#  
���0 c                   �  ���  ���1 0 PreB  ���        �  [���6  O���  m���>  [��� PreC    �6  O���(  O���1 f                  �6  [���(  [���0 g                   �  U���  U���1 0 PreC  m���        �V  ����b  ����l  �����  ���� CirALL    �V  ����V  ����1 [                  �b  ����b  ����0 \                   �\  ����\  ����1 0 CirALLl  ����        ��  �����  �����  �����  ����  Z     ��  �����  ����1 1 Z�  ����          ��  Cnand3�   `���   <���                       ��   Z����   Z���1 1                  ��   N����   N���1 1                  ��   B����   B���0 0                   �  N���  N���1 1                  ��  Cnand2�   *���  ���                       ��   ����   ���1 1                  ��   ����   ���1 1                   �  ����   ���0 0                  <�j  E����  !���                       �j  9���x  9���1 1                  �j  -���x  -���0 0                   ��  3����  3���1 1                  �C   ����s   ����P   ����f   ���� X     �C   ����Q   ����1 #                  �C   ����Q   ����0 $                   �s   ����e   ����1 0 Xs   ����        ��  Cnor3p  �����  ����                       �p  �����  ����1 1                  �p  �����  ����1 1                  �p  �����  ����1 1                   ��  �����  ����0 0                  �� 	 Cinverter`   	����   ����                      �r   	���r   ����1 1                   �r   ����r   ����0 0                  6��  ����  ����                       ��  �����  ����1 1                  ��  �����  ����1 1                  ��  �����  ����1 1                   �   �����  ����0 0                  <�8  �����  g���                       �8  ���F  ���0 0                  �8  s���F  s���1 1                   ��  y���t  y���1 1                  <��  h����  D���                       ��  \����  \���0 0                  ��  P����  P���1 1                   ��  V����  V���1 1                   ��  Cnet1  ��  Csegment[  ����[  ���b�[  ����[  ����b�[  ����  ���b��  ����  ���b��  ����  ���b�[  Q����  Q���b�[  ����[  Q���b��  Q����  Q���b�[  �����  ����b�[  Q���[  ����b��  �����  ����     # `�0  b�`  ����`  i���b�  i���`  i���b�  i���  i���b�`  ����`  ����    `�0  b�g  ����g  ����b�  ����g  ����b�  ����  ����b�g  ����g  ����    `�1  b��  �����  ����b�  �����  ����b�  ����  ����b��  �����  ����   ' `�1  b��  �����  ���b�  ����  ���b�  ���  ���b��  �����  ����   + `�1  b��  Z����  U���b�  U����  U���b�  U���  U���b��  Z����  Z���   / `�1  b��  �����  ����b�E  �����  ����b�\  ����\  ����b��  �����  ����b�E  ����E  +���b��  +���E  +���b��  +����  +���b�E  �����  ����b�E  ����E  ����b��  �����  ����b�E  ����E  ����b�\  ����E  ����     3 `�0 	 b�  ���  ����b�A  ����  ����b�  ���  ���b�A  ����A  i���b��  i���A  i���b��  i����  i���b�A  �����   ����b��   �����   B���b��   B����   B���  :   `�1  b��   ���s   ���b�s   ����s   ���b�s   ����s   ����b��   ����   ���b��   ����   ���b��   ����   ����b��  �����   ����b�s   ���r   ���b�r   ���r   	���b�r   	���r   	���b��  �����  ���� > Q T  H `�1  b�j  9���  9���b�  N���  9���b�  N���  N���b�j  9���j  9��� B  ; `�0  b�j  -���  -���b�  ���  -���b�  ���  ���b�j  -���j  -��� C  @ `�1  b��  4����  4���b��  3����  4���b��  3����  3���b��  4����  4���   D `�1  b�  Q���   ���b�   ���   ���b�  Q���  Q���b�  ����  ����b�4  ����p  ����b�p  ����p  ����b�   ���  ����b�  �����   ����b��   Z����   ����b��   Z����   Z���b�  ����4  ����b�4  ����4  ����b��  ����4  ����b��  �����  ���� K 8 U   `�0  b��  �����  ����b��  �����  ����b��  �����  ����b��  �����  ����   N `�1  b�  ����  ����b�f  ����  ����b�  ����  ����b�p  ����p  ����b�f  �����   ����b��   �����   N���b��   N����   N���b��   N����   N���b�f  ����p  ����b�f  ����f  ����b�f  ����f  ����b�f  �����  ����b��  �����  ���� L 9 V   `�1  b�|  4���*  4���b�  4���  4���b�|  E���|  E���b�  4���*  4���b�*  4���*  ����b�O  ����*  ����b��   �����   ���b��   ����   ���b��   ����   ���b��   ����O  ����b�O  ����O  ����b�p  ����O  ����b�p  ����p  ����b�|  E���|  4���b�O  ����O  L���b�O  L����  L���b��  P����  L���b��  P����  P���b��  P����  P���b��  P����  P���  ? M ^   `�1  b��  y����  y���b��  �����  y���b��  �����  ����b��  y����  y��� 5  [ `�0  b��  \���r   \���b�r   ����r   \���b�r   ����r   ����b��  \����  \��� ]  R `�0  b�8  ���   ���b�   ����   ���b�   ����   ����b�8  ���8  ��� Y  W `�1  b�8  s����  s���b��  V����  s���b��  V����  V���b�8  s���8  s��� Z  _   joshua